`timescale 1ns/1ps
`include "verilog_spice/cod_decod.v"
module cod_decod_tb;
    initial begin
        
    end
endmodule