module encoder;
    
endmodule